
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity tb_sobelProc is
end entity tb_sobelProc;

architecture archi_tb_sobelProc of tb_sobelProc is
  component sobelProc is
    Port ( clk,reset		: in STD_LOGIC;
		   I_go	   			: in STD_LOGIC;
		   -- interface avec la mémoire IN (lecture)
		   O_enM_R		 	: out STD_LOGIC;
		   O_ADR_R		 	: out STD_LOGIC_VECTOR (13 downto 0); 
		   I_pixel 			: in  STD_LOGIC_VECTOR (7 downto 0); -- Pixel from memory IN
		   -- interface avec la mémoire OUT (écriture)
		   O_enM_W		 	: out STD_LOGIC;		   
		   O_ADR_W	 	 	: out STD_LOGIC_VECTOR (13 downto 0); 
		   O_pixEdge 		: out  STD_LOGIC; -- Edge to memory OUT
		   -- signal de commande vers le contrôleur VGA		   		   
		   O_StartDisplay	: out STD_LOGIC
		   ); 
  end component sobelProc;

signal S_clk             :  STD_LOGIC := '0';
signal S_reset	       :  STD_LOGIC;
signal S_go	   		   :  STD_LOGIC;
signal S_enM_R		   :  STD_LOGIC;
signal S_ADR_R		   :  STD_LOGIC_VECTOR (13 downto 0);
signal S_pixel 		   :  STD_LOGIC_VECTOR (7 downto 0);
signal S_enM_W		   :  STD_LOGIC;
signal S_ADR_W	 	   :  STD_LOGIC_VECTOR (13 downto 0);
signal S_pixEdge 	   :  STD_LOGIC;
signal S_StartDisplay  :  STD_LOGIC;
  


begin
  S_pixel <= "00000111" after 0 ns, "11111111" after 10 ns, "01100111" after 20 ns, "01111011" after 30 ns, "00000111" after 40 ns, "11111111" after 50 ns, "01100111" after 60 ns, "01111011" after 70 ns, "00000111" after 80 ns, "11111111" after 90 ns, "01100111" after 100 ns, "01111011" after 110 ns, "00000111" after 120 ns, "11111111" after 130 ns, "01100111" after 140 ns, "01111011" after 150 ns, "00000111" after 160 ns, "11111111" after 170 ns, "01100111" after 180 ns, "01111011" after 190 ns, "00000111" after 200 ns, "11111111" after 210 ns, "01100111" after 220 ns, "01111011" after 230 ns, "00000111" after 240 ns, "11111111" after 250 ns, "01100111" after 260 ns, "01111011" after 270 ns, "00000111" after 280 ns, "11111111" after 290 ns, "01100111" after 300 ns, "01111011" after 310 ns, "00000111" after 320 ns, "11111111" after 330 ns, "01100111" after 340 ns, "01111011" after 350 ns, "00000111" after 360 ns, "11111111" after 370 ns, "01100111" after 380 ns, "01111011" after 390 ns, "00000111" after 400 ns, "11111111" after 410 ns, "01100111" after 420 ns, "01111011" after 430 ns, "00000111" after 440 ns, "11111111" after 450 ns, "01100111" after 460 ns, "01111011" after 470 ns, "00000111" after 480 ns, "11111111" after 490 ns, "01100111" after 500 ns, "01111011" after 510 ns, "00000111" after 520 ns, "11111111" after 530 ns, "01100111" after 540 ns, "01111011" after 550 ns, "00000111" after 560 ns, "11111111" after 570 ns, "01100111" after 580 ns, "01111011" after 590 ns, "00000111" after 600 ns, "11111111" after 610 ns, "01100111" after 620 ns, "01111011" after 630 ns, "00000111" after 640 ns, "11111111" after 650 ns, "01100111" after 660 ns, "01111011" after 670 ns, "00000111" after 680 ns, "11111111" after 690 ns, "01100111" after 700 ns, "01111011" after 710 ns, "00000111" after 720 ns, "11111111" after 730 ns, "01100111" after 740 ns, "01111011" after 750 ns, "00000111" after 760 ns, "11111111" after 770 ns, "01100111" after 780 ns, "01111011" after 790 ns, "00000111" after 800 ns, "11111111" after 810 ns, "01100111" after 820 ns, "01111011" after 830 ns, "00000111" after 840 ns, "11111111" after 850 ns, "01100111" after 860 ns, "01111011" after 870 ns, "00000111" after 880 ns, "11111111" after 890 ns, "01100111" after 900 ns, "01111011" after 910 ns, "00000111" after 920 ns, "11111111" after 930 ns, "01100111" after 940 ns, "01111011" after 950 ns, "00000111" after 960 ns, "11111111" after 970 ns, "01100111" after 980 ns, "01111011" after 990 ns, "00000111" after 1000 ns, "11111111" after 1010 ns, "01100111" after 1020 ns, "01111011" after 1030 ns, "00000111" after 1040 ns, "11111111" after 1050 ns, "01100111" after 1060 ns, "01111011" after 1070 ns, "00000111" after 1080 ns, "11111111" after 1090 ns, "01100111" after 1100 ns, "01111011" after 1110 ns, "00000111" after 1120 ns, "11111111" after 1130 ns, "01100111" after 1140 ns, "01111011" after 1150 ns, "00000111" after 1160 ns, "11111111" after 1170 ns, "01100111" after 1180 ns, "01111011" after 1190 ns, "00000111" after 1200 ns, "11111111" after 1210 ns, "01100111" after 1220 ns, "01111011" after 1230 ns, "00000111" after 1240 ns, "11111111" after 1250 ns, "01100111" after 1260 ns, "01111011" after 1270 ns, "00000111" after 1280 ns, "11111111" after 1290 ns, "01100111" after 1300 ns, "01111011" after 1310 ns, "00000111" after 1320 ns, "11111111" after 1330 ns, "01100111" after 1340 ns, "01111011" after 1350 ns, "00000111" after 1360 ns, "11111111" after 1370 ns, "01100111" after 1380 ns, "01111011" after 1390 ns, "00000111" after 1400 ns, "11111111" after 1410 ns, "01100111" after 1420 ns, "01111011" after 1430 ns, "00000111" after 1440 ns, "11111111" after 1450 ns, "01100111" after 1460 ns, "01111011" after 1470 ns, "00000111" after 1480 ns, "11111111" after 1490 ns, "01100111" after 1500 ns, "01111011" after 1510 ns, "00000111" after 1520 ns, "11111111" after 1530 ns, "01100111" after 1540 ns, "01111011" after 1550 ns, "00000111" after 1560 ns, "11111111" after 1570 ns, "01100111" after 1580 ns, "01111011" after 1590 ns, "00000111" after 1600 ns, "11111111" after 1610 ns, "01100111" after 1620 ns, "01111011" after 1630 ns, "00000111" after 1640 ns, "11111111" after 1650 ns, "01100111" after 1660 ns, "01111011" after 1670 ns, "00000111" after 1680 ns, "11111111" after 1690 ns, "01100111" after 1700 ns, "01111011" after 1710 ns, "00000111" after 1720 ns, "11111111" after 1730 ns, "01100111" after 1740 ns, "01111011" after 1750 ns, "00000111" after 1760 ns, "11111111" after 1770 ns, "01100111" after 1780 ns, "01111011" after 1790 ns, "00000111" after 1800 ns, "11111111" after 1810 ns, "01100111" after 1820 ns, "01111011" after 1830 ns, "00000111" after 1840 ns, "11111111" after 1850 ns, "01100111" after 1860 ns, "01111011" after 1870 ns, "00000111" after 1880 ns, "11111111" after 1890 ns, "01100111" after 1900 ns, "01111011" after 1910 ns, "00000111" after 1920 ns, "11111111" after 1930 ns, "01100111" after 1940 ns, "01111011" after 1950 ns, "00000111" after 1960 ns, "11111111" after 1970 ns, "01100111" after 1980 ns, "01111011" after 1990 ns, "00000111" after 2000 ns, "11111111" after 2010 ns, "01100111" after 2020 ns, "01111011" after 2030 ns, "00000111" after 2040 ns, "11111111" after 2050 ns, "01100111" after 2060 ns, "01111011" after 2070 ns, "00000111" after 2080 ns, "11111111" after 2090 ns, "01100111" after 2100 ns, "01111011" after 2110 ns, "00000111" after 2120 ns, "11111111" after 2130 ns, "01100111" after 2140 ns, "01111011" after 2150 ns, "00000111" after 2160 ns, "11111111" after 2170 ns, "01100111" after 2180 ns, "01111011" after 2190 ns, "00000111" after 2200 ns, "11111111" after 2210 ns, "01100111" after 2220 ns, "01111011" after 2230 ns, "00000111" after 2240 ns, "11111111" after 2250 ns, "01100111" after 2260 ns, "01111011" after 2270 ns, "00000111" after 2280 ns, "11111111" after 2290 ns, "01100111" after 2300 ns, "01111011" after 2310 ns, "00000111" after 2320 ns, "11111111" after 2330 ns, "01100111" after 2340 ns, "01111011" after 2350 ns, "00000111" after 2360 ns, "11111111" after 2370 ns, "01100111" after 2380 ns, "01111011" after 2390 ns, "00000111" after 2400 ns, "11111111" after 2410 ns, "01100111" after 2420 ns, "01111011" after 2430 ns, "00000111" after 2440 ns, "11111111" after 2450 ns, "01100111" after 2460 ns, "01111011" after 2470 ns, "00000111" after 2480 ns, "11111111" after 2490 ns, "01100111" after 2500 ns, "01111011" after 2510 ns, "00000111" after 2520 ns, "11111111" after 2530 ns, "01100111" after 2540 ns, "01111011" after 2550 ns, "00000111" after 2560 ns, "11111111" after 2570 ns, "01100111" after 2580 ns, "01111011" after 2590 ns, "00000111" after 2600 ns, "11111111" after 2610 ns, "01100111" after 2620 ns, "01111011" after 2630 ns, "00000111" after 2640 ns, "11111111" after 2650 ns, "01100111" after 2660 ns, "01111011" after 2670 ns, "00000111" after 2680 ns, "11111111" after 2690 ns, "01100111" after 2700 ns, "01111011" after 2710 ns, "00000111" after 2720 ns, "11111111" after 2730 ns, "01100111" after 2740 ns, "01111011" after 2750 ns, "00000111" after 2760 ns, "11111111" after 2770 ns, "01100111" after 2780 ns, "01111011" after 2790 ns, "00000111" after 2800 ns, "11111111" after 2810 ns, "01100111" after 2820 ns, "01111011" after 2830 ns, "00000111" after 2840 ns, "11111111" after 2850 ns, "01100111" after 2860 ns, "01111011" after 2870 ns, "00000111" after 2880 ns, "11111111" after 2890 ns, "01100111" after 2900 ns, "01111011" after 2910 ns, "00000111" after 2920 ns, "11111111" after 2930 ns, "01100111" after 2940 ns, "01111011" after 2950 ns, "00000111" after 2960 ns, "11111111" after 2970 ns, "01100111" after 2980 ns, "01111011" after 2990 ns, "00000111" after 3000 ns, "11111111" after 3010 ns, "01100111" after 3020 ns, "01111011" after 3030 ns, "00000111" after 3040 ns, "11111111" after 3050 ns, "01100111" after 3060 ns, "01111011" after 3070 ns, "00000111" after 3080 ns, "11111111" after 3090 ns, "01100111" after 3100 ns, "01111011" after 3110 ns, "00000111" after 3120 ns, "11111111" after 3130 ns, "01100111" after 3140 ns, "01111011" after 3150 ns, "00000111" after 3160 ns, "11111111" after 3170 ns, "01100111" after 3180 ns, "01111011" after 3190 ns, "00000111" after 3200 ns, "11111111" after 3210 ns, "01100111" after 3220 ns, "01111011" after 3230 ns, "00000111" after 3240 ns, "11111111" after 3250 ns, "01100111" after 3260 ns, "01111011" after 3270 ns, "00000111" after 3280 ns, "11111111" after 3290 ns, "01100111" after 3300 ns, "01111011" after 3310 ns, "00000111" after 3320 ns, "11111111" after 3330 ns, "01100111" after 3340 ns, "01111011" after 3350 ns, "00000111" after 3360 ns, "11111111" after 3370 ns, "01100111" after 3380 ns, "01111011" after 3390 ns, "00000111" after 3400 ns, "11111111" after 3410 ns, "01100111" after 3420 ns, "01111011" after 3430 ns, "00000111" after 3440 ns, "11111111" after 3450 ns, "01100111" after 3460 ns, "01111011" after 3470 ns, "00000111" after 3480 ns, "11111111" after 3490 ns, "01100111" after 3500 ns, "01111011" after 3510 ns, "00000111" after 3520 ns, "11111111" after 3530 ns, "01100111" after 3540 ns, "01111011" after 3550 ns, "00000111" after 3560 ns, "11111111" after 3570 ns, "01100111" after 3580 ns, "01111011" after 3590 ns, "00000111" after 3600 ns, "11111111" after 3610 ns, "01100111" after 3620 ns, "01111011" after 3630 ns, "00000111" after 3640 ns, "11111111" after 3650 ns, "01100111" after 3660 ns, "01111011" after 3670 ns, "00000111" after 3680 ns, "11111111" after 3690 ns, "01100111" after 3700 ns, "01111011" after 3710 ns, "00000111" after 3720 ns, "11111111" after 3730 ns, "01100111" after 3740 ns, "01111011" after 3750 ns, "00000111" after 3760 ns, "11111111" after 3770 ns, "01100111" after 3780 ns, "01111011" after 3790 ns, "00000111" after 3800 ns, "11111111" after 3810 ns, "01100111" after 3820 ns, "01111011" after 3830 ns, "00000111" after 3840 ns, "11111111" after 3850 ns, "01100111" after 3860 ns, "01111011" after 3870 ns, "00000111" after 3880 ns, "11111111" after 3890 ns, "01100111" after 3900 ns, "01111011" after 3910 ns, "00000111" after 3920 ns, "11111111" after 3930 ns, "01100111" after 3940 ns, "01111011" after 3950 ns, "00000111" after 3960 ns, "11111111" after 3970 ns, "01100111" after 3980 ns, "01111011" after 3990 ns, "00000111" after 4000 ns, "11111111" after 4010 ns, "01100111" after 4020 ns, "01111011" after 4030 ns, "00000111" after 4040 ns, "11111111" after 4050 ns, "01100111" after 4060 ns, "01111011" after 4070 ns, "00000111" after 4080 ns, "11111111" after 4090 ns, "01100111" after 4100 ns, "01111011" after 4110 ns, "00000111" after 4120 ns, "11111111" after 4130 ns, "01100111" after 4140 ns, "01111011" after 4150 ns, "00000111" after 4160 ns, "11111111" after 4170 ns, "01100111" after 4180 ns, "01111011" after 4190 ns, "00000111" after 4200 ns, "11111111" after 4210 ns, "01100111" after 4220 ns, "01111011" after 4230 ns, "00000111" after 4240 ns, "11111111" after 4250 ns, "01100111" after 4260 ns, "01111011" after 4270 ns, "00000111" after 4280 ns, "11111111" after 4290 ns, "01100111" after 4300 ns, "01111011" after 4310 ns, "00000111" after 4320 ns, "11111111" after 4330 ns, "01100111" after 4340 ns, "01111011" after 4350 ns, "00000111" after 4360 ns, "11111111" after 4370 ns, "01100111" after 4380 ns, "01111011" after 4390 ns, "00000111" after 4400 ns, "11111111" after 4410 ns, "01100111" after 4420 ns, "01111011" after 4430 ns, "00000111" after 4440 ns, "11111111" after 4450 ns, "01100111" after 4460 ns, "01111011" after 4470 ns, "00000111" after 4480 ns, "11111111" after 4490 ns, "01100111" after 4500 ns, "01111011" after 4510 ns, "00000111" after 4520 ns, "11111111" after 4530 ns, "01100111" after 4540 ns, "01111011" after 4550 ns, "00000111" after 4560 ns, "11111111" after 4570 ns, "01100111" after 4580 ns, "01111011" after 4590 ns, "00000111" after 4600 ns, "11111111" after 4610 ns, "01100111" after 4620 ns, "01111011" after 4630 ns, "00000111" after 4640 ns, "11111111" after 4650 ns, "01100111" after 4660 ns, "01111011" after 4670 ns, "00000111" after 4680 ns, "11111111" after 4690 ns, "01100111" after 4700 ns, "01111011" after 4710 ns, "00000111" after 4720 ns, "11111111" after 4730 ns, "01100111" after 4740 ns, "01111011" after 4750 ns, "00000111" after 4760 ns, "11111111" after 4770 ns, "01100111" after 4780 ns, "01111011" after 4790 ns, "00000111" after 4800 ns, "11111111" after 4810 ns, "01100111" after 4820 ns, "01111011" after 4830 ns, "00000111" after 4840 ns, "11111111" after 4850 ns, "01100111" after 4860 ns, "01111011" after 4870 ns, "00000111" after 4880 ns, "11111111" after 4890 ns, "01100111" after 4900 ns, "01111011" after 4910 ns, "00000111" after 4920 ns, "11111111" after 4930 ns, "01100111" after 4940 ns, "01111011" after 4950 ns, "00000111" after 4960 ns, "11111111" after 4970 ns, "01100111" after 4980 ns, "01111011" after 4990 ns, "00000111" after 5000 ns, "11111111" after 5010 ns, "01100111" after 5020 ns, "01111011" after 5030 ns, "00000111" after 5040 ns, "11111111" after 5050 ns, "01100111" after 5060 ns, "01111011" after 5070 ns, "00000111" after 5080 ns, "11111111" after 5090 ns, "01100111" after 5100 ns, "01111011" after 5110 ns, "00000111" after 5120 ns, "11111111" after 5130 ns, "01100111" after 5140 ns, "01111011" after 5150 ns, "00000111" after 5160 ns, "11111111" after 5170 ns, "01100111" after 5180 ns, "01111011" after 5190 ns, "00000111" after 5200 ns, "11111111" after 5210 ns, "01100111" after 5220 ns, "01111011" after 5230 ns, "00000111" after 5240 ns, "11111111" after 5250 ns, "01100111" after 5260 ns, "01111011" after 5270 ns, "00000111" after 5280 ns, "11111111" after 5290 ns, "01100111" after 5300 ns, "01111011" after 5310 ns, "00000111" after 5320 ns, "11111111" after 5330 ns, "01100111" after 5340 ns, "01111011" after 5350 ns, "00000111" after 5360 ns, "11111111" after 5370 ns, "01100111" after 5380 ns, "01111011" after 5390 ns, "00000111" after 5400 ns, "11111111" after 5410 ns, "01100111" after 5420 ns, "01111011" after 5430 ns, "00000111" after 5440 ns, "11111111" after 5450 ns, "01100111" after 5460 ns, "01111011" after 5470 ns, "00000111" after 5480 ns, "11111111" after 5490 ns, "01100111" after 5500 ns, "01111011" after 5510 ns, "00000111" after 5520 ns, "11111111" after 5530 ns, "01100111" after 5540 ns, "01111011" after 5550 ns, "00000111" after 5560 ns, "11111111" after 5570 ns, "01100111" after 5580 ns, "01111011" after 5590 ns, "00000111" after 5600 ns, "11111111" after 5610 ns, "01100111" after 5620 ns, "01111011" after 5630 ns, "00000111" after 5640 ns, "11111111" after 5650 ns, "01100111" after 5660 ns, "01111011" after 5670 ns, "00000111" after 5680 ns, "11111111" after 5690 ns, "01100111" after 5700 ns, "01111011" after 5710 ns, "00000111" after 5720 ns, "11111111" after 5730 ns, "01100111" after 5740 ns, "01111011" after 5750 ns, "00000111" after 5760 ns, "11111111" after 5770 ns, "01100111" after 5780 ns, "01111011" after 5790 ns, "00000111" after 5800 ns, "11111111" after 5810 ns, "01100111" after 5820 ns, "01111011" after 5830 ns, "00000111" after 5840 ns, "11111111" after 5850 ns, "01100111" after 5860 ns, "01111011" after 5870 ns, "00000111" after 5880 ns, "11111111" after 5890 ns, "01100111" after 5900 ns, "01111011" after 5910 ns, "00000111" after 5920 ns, "11111111" after 5930 ns, "01100111" after 5940 ns, "01111011" after 5950 ns, "00000111" after 5960 ns, "11111111" after 5970 ns, "01100111" after 5980 ns, "01111011" after 5990 ns, "00000111" after 6000 ns, "11111111" after 6010 ns, "01100111" after 6020 ns, "01111011" after 6030 ns, "00000111" after 6040 ns, "11111111" after 6050 ns, "01100111" after 6060 ns, "01111011" after 6070 ns, "00000111" after 6080 ns, "11111111" after 6090 ns, "01100111" after 6100 ns, "01111011" after 6110 ns, "00000111" after 6120 ns, "11111111" after 6130 ns, "01100111" after 6140 ns, "01111011" after 6150 ns, "00000111" after 6160 ns, "11111111" after 6170 ns, "01100111" after 6180 ns, "01111011" after 6190 ns, "00000111" after 6200 ns, "11111111" after 6210 ns, "01100111" after 6220 ns, "01111011" after 6230 ns, "00000111" after 6240 ns, "11111111" after 6250 ns, "01100111" after 6260 ns, "01111011" after 6270 ns, "00000111" after 6280 ns, "11111111" after 6290 ns, "01100111" after 6300 ns, "01111011" after 6310 ns, "00000111" after 6320 ns, "11111111" after 6330 ns, "01100111" after 6340 ns, "01111011" after 6350 ns, "00000111" after 6360 ns, "11111111" after 6370 ns, "01100111" after 6380 ns, "01111011" after 6390 ns, "00000111" after 6400 ns, "11111111" after 6410 ns, "01100111" after 6420 ns, "01111011" after 6430 ns, "00000111" after 6440 ns, "11111111" after 6450 ns, "01100111" after 6460 ns, "01111011" after 6470 ns, "00000111" after 6480 ns, "11111111" after 6490 ns, "01100111" after 6500 ns, "01111011" after 6510 ns, "00000111" after 6520 ns, "11111111" after 6530 ns, "01100111" after 6540 ns, "01111011" after 6550 ns, "00000111" after 6560 ns, "11111111" after 6570 ns, "01100111" after 6580 ns, "01111011" after 6590 ns, "00000111" after 6600 ns, "11111111" after 6610 ns, "01100111" after 6620 ns, "01111011" after 6630 ns, "00000111" after 6640 ns, "11111111" after 6650 ns, "01100111" after 6660 ns, "01111011" after 6670 ns, "00000111" after 6680 ns, "11111111" after 6690 ns, "01100111" after 6700 ns, "01111011" after 6710 ns, "00000111" after 6720 ns, "11111111" after 6730 ns, "01100111" after 6740 ns, "01111011" after 6750 ns, "00000111" after 6760 ns, "11111111" after 6770 ns, "01100111" after 6780 ns, "01111011" after 6790 ns, "00000111" after 6800 ns, "11111111" after 6810 ns, "01100111" after 6820 ns, "01111011" after 6830 ns, "00000111" after 6840 ns, "11111111" after 6850 ns, "01100111" after 6860 ns, "01111011" after 6870 ns, "00000111" after 6880 ns, "11111111" after 6890 ns, "01100111" after 6900 ns, "01111011" after 6910 ns, "00000111" after 6920 ns, "11111111" after 6930 ns, "01100111" after 6940 ns, "01111011" after 6950 ns, "00000111" after 6960 ns, "11111111" after 6970 ns, "01100111" after 6980 ns, "01111011" after 6990 ns, "00000111" after 7000 ns, "11111111" after 7010 ns, "01100111" after 7020 ns, "01111011" after 7030 ns, "00000111" after 7040 ns, "11111111" after 7050 ns, "01100111" after 7060 ns, "01111011" after 7070 ns, "00000111" after 7080 ns, "11111111" after 7090 ns, "01100111" after 7100 ns, "01111011" after 7110 ns, "00000111" after 7120 ns, "11111111" after 7130 ns, "01100111" after 7140 ns, "01111011" after 7150 ns, "00000111" after 7160 ns, "11111111" after 7170 ns, "01100111" after 7180 ns, "01111011" after 7190 ns, "00000111" after 7200 ns, "11111111" after 7210 ns, "01100111" after 7220 ns, "01111011" after 7230 ns, "00000111" after 7240 ns, "11111111" after 7250 ns, "01100111" after 7260 ns, "01111011" after 7270 ns, "00000111" after 7280 ns, "11111111" after 7290 ns, "01100111" after 7300 ns, "01111011" after 7310 ns, "00000111" after 7320 ns, "11111111" after 7330 ns, "01100111" after 7340 ns, "01111011" after 7350 ns, "00000111" after 7360 ns, "11111111" after 7370 ns, "01100111" after 7380 ns, "01111011" after 7390 ns, "00000111" after 7400 ns, "11111111" after 7410 ns, "01100111" after 7420 ns, "01111011" after 7430 ns, "00000111" after 7440 ns, "11111111" after 7450 ns, "01100111" after 7460 ns, "01111011" after 7470 ns, "00000111" after 7480 ns, "11111111" after 7490 ns, "01100111" after 7500 ns, "01111011" after 7510 ns, "00000111" after 7520 ns, "11111111" after 7530 ns, "01100111" after 7540 ns, "01111011" after 7550 ns, "00000111" after 7560 ns, "11111111" after 7570 ns, "01100111" after 7580 ns, "01111011" after 7590 ns, "00000111" after 7600 ns, "11111111" after 7610 ns, "01100111" after 7620 ns, "01111011" after 7630 ns, "00000111" after 7640 ns, "11111111" after 7650 ns, "01100111" after 7660 ns, "01111011" after 7670 ns, "00000111" after 7680 ns, "11111111" after 7690 ns, "01100111" after 7700 ns, "01111011" after 7710 ns, "00000111" after 7720 ns, "11111111" after 7730 ns, "01100111" after 7740 ns, "01111011" after 7750 ns, "00000111" after 7760 ns, "11111111" after 7770 ns, "01100111" after 7780 ns, "01111011" after 7790 ns, "00000111" after 7800 ns, "11111111" after 7810 ns, "01100111" after 7820 ns, "01111011" after 7830 ns, "00000111" after 7840 ns, "11111111" after 7850 ns, "01100111" after 7860 ns, "01111011" after 7870 ns, "00000111" after 7880 ns, "11111111" after 7890 ns, "01100111" after 7900 ns, "01111011" after 7910 ns, "00000111" after 7920 ns, "11111111" after 7930 ns, "01100111" after 7940 ns, "01111011" after 7950 ns, "00000111" after 7960 ns, "11111111" after 7970 ns, "01100111" after 7980 ns, "01111011" after 7990 ns, "00000111" after 8000 ns, "11111111" after 8010 ns, "01100111" after 8020 ns, "01111011" after 8030 ns, "00000111" after 8040 ns, "11111111" after 8050 ns, "01100111" after 8060 ns, "01111011" after 8070 ns, "00000111" after 8080 ns, "11111111" after 8090 ns, "01100111" after 8100 ns, "01111011" after 8110 ns, "00000111" after 8120 ns, "11111111" after 8130 ns, "01100111" after 8140 ns, "01111011" after 8150 ns, "00000111" after 8160 ns, "11111111" after 8170 ns, "01100111" after 8180 ns, "01111011" after 8190 ns, "00000111" after 8200 ns, "11111111" after 8210 ns, "01100111" after 8220 ns, "01111011" after 8230 ns, "00000111" after 8240 ns, "11111111" after 8250 ns, "01100111" after 8260 ns, "01111011" after 8270 ns, "00000111" after 8280 ns, "11111111" after 8290 ns, "01100111" after 8300 ns, "01111011" after 8310 ns, "00000111" after 8320 ns, "11111111" after 8330 ns, "01100111" after 8340 ns, "01111011" after 8350 ns, "00000111" after 8360 ns, "11111111" after 8370 ns, "01100111" after 8380 ns, "01111011" after 8390 ns, "00000111" after 8400 ns, "11111111" after 8410 ns, "01100111" after 8420 ns, "01111011" after 8430 ns, "00000111" after 8440 ns, "11111111" after 8450 ns, "01100111" after 8460 ns, "01111011" after 8470 ns, "00000111" after 8480 ns, "11111111" after 8490 ns, "01100111" after 8500 ns, "01111011" after 8510 ns, "00000111" after 8520 ns, "11111111" after 8530 ns, "01100111" after 8540 ns, "01111011" after 8550 ns, "00000111" after 8560 ns, "11111111" after 8570 ns, "01100111" after 8580 ns, "01111011" after 8590 ns, "00000111" after 8600 ns, "11111111" after 8610 ns, "01100111" after 8620 ns, "01111011" after 8630 ns, "00000111" after 8640 ns, "11111111" after 8650 ns, "01100111" after 8660 ns, "01111011" after 8670 ns, "00000111" after 8680 ns, "11111111" after 8690 ns, "01100111" after 8700 ns, "01111011" after 8710 ns, "00000111" after 8720 ns, "11111111" after 8730 ns, "01100111" after 8740 ns, "01111011" after 8750 ns, "00000111" after 8760 ns, "11111111" after 8770 ns, "01100111" after 8780 ns, "01111011" after 8790 ns, "00000111" after 8800 ns, "11111111" after 8810 ns, "01100111" after 8820 ns, "01111011" after 8830 ns, "00000111" after 8840 ns, "11111111" after 8850 ns, "01100111" after 8860 ns, "01111011" after 8870 ns, "00000111" after 8880 ns, "11111111" after 8890 ns, "01100111" after 8900 ns, "01111011" after 8910 ns, "00000111" after 8920 ns, "11111111" after 8930 ns, "01100111" after 8940 ns, "01111011" after 8950 ns, "00000111" after 8960 ns, "11111111" after 8970 ns, "01100111" after 8980 ns, "01111011" after 8990 ns, "00000111" after 9000 ns, "11111111" after 9010 ns, "01100111" after 9020 ns, "01111011" after 9030 ns, "00000111" after 9040 ns, "11111111" after 9050 ns, "01100111" after 9060 ns, "01111011" after 9070 ns, "00000111" after 9080 ns, "11111111" after 9090 ns, "01100111" after 9100 ns, "01111011" after 9110 ns, "00000111" after 9120 ns, "11111111" after 9130 ns, "01100111" after 9140 ns, "01111011" after 9150 ns, "00000111" after 9160 ns, "11111111" after 9170 ns, "01100111" after 9180 ns, "01111011" after 9190 ns, "00000111" after 9200 ns, "11111111" after 9210 ns, "01100111" after 9220 ns, "01111011" after 9230 ns, "00000111" after 9240 ns, "11111111" after 9250 ns, "01100111" after 9260 ns, "01111011" after 9270 ns, "00000111" after 9280 ns, "11111111" after 9290 ns, "01100111" after 9300 ns, "01111011" after 9310 ns, "00000111" after 9320 ns, "11111111" after 9330 ns, "01100111" after 9340 ns, "01111011" after 9350 ns, "00000111" after 9360 ns, "11111111" after 9370 ns, "01100111" after 9380 ns, "01111011" after 9390 ns, "00000111" after 9400 ns, "11111111" after 9410 ns, "01100111" after 9420 ns, "01111011" after 9430 ns, "00000111" after 9440 ns, "11111111" after 9450 ns, "01100111" after 9460 ns, "01111011" after 9470 ns, "00000111" after 9480 ns, "11111111" after 9490 ns, "01100111" after 9500 ns, "01111011" after 9510 ns, "00000111" after 9520 ns, "11111111" after 9530 ns, "01100111" after 9540 ns, "01111011" after 9550 ns, "00000111" after 9560 ns, "11111111" after 9570 ns, "01100111" after 9580 ns, "01111011" after 9590 ns, "00000111" after 9600 ns, "11111111" after 9610 ns, "01100111" after 9620 ns, "01111011" after 9630 ns, "00000111" after 9640 ns, "11111111" after 9650 ns, "01100111" after 9660 ns, "01111011" after 9670 ns, "00000111" after 9680 ns, "11111111" after 9690 ns, "01100111" after 9700 ns, "01111011" after 9710 ns, "00000111" after 9720 ns, "11111111" after 9730 ns, "01100111" after 9740 ns, "01111011" after 9750 ns, "00000111" after 9760 ns, "11111111" after 9770 ns, "01100111" after 9780 ns, "01111011" after 9790 ns, "00000111" after 9800 ns, "11111111" after 9810 ns, "01100111" after 9820 ns, "01111011" after 9830 ns, "00000111" after 9840 ns, "11111111" after 9850 ns, "01100111" after 9860 ns, "01111011" after 9870 ns, "00000111" after 9880 ns, "11111111" after 9890 ns, "01100111" after 9900 ns, "01111011" after 9910 ns, "00000111" after 9920 ns, "11111111" after 9930 ns, "01100111" after 9940 ns, "01111011" after 9950 ns, "00000111" after 9960 ns, "11111111" after 9970 ns, "01100111" after 9980 ns, "01111011" after 9990 ns;

  
  S_clk <= not S_clk after 5 ns;
  S_reset <= '1', '0' after 64 ns;
  S_go <= '0', '1' after 164 ns, '0' after 264 ns;  

  sobelProc_1 : entity work.sobelProc
    port map (
      clk               => S_clk          ,
      reset	            => S_reset	      ,
      I_go	   		    => S_go	   		  ,
      O_enM_R		    => S_enM_R		  ,
      O_ADR_R		    => S_ADR_R		  ,
      I_pixel 		    => S_pixel 		  ,
      O_enM_W		    => S_enM_W		  ,
      O_ADR_W	 	    => S_ADR_W	 	  ,
      O_pixEdge 	    => S_pixEdge 	  ,
      O_StartDisplay    => S_StartDisplay 
	  );
      

end architecture archi_tb_sobelProc;
